module ADDER (
	input [7:0] a,
	input [7:0] b,
	output [8:0] do,
	);

assign do = a + b;

endmodule
